interface adder_intf (input clk, rst);
  
endinterface