interface adder_intf (input clk, rst);
  bit a;
  bit b;
  bit c;
  bit sum;
  bit carry;
endinterface