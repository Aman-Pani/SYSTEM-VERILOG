// https://www.edaplayground.com/x/Hf85

// parameterized_class  :  
// scope resolution     :  
// casting              :
