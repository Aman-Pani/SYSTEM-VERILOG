// `include "randomization_01.sv"
// `include "constraint_inside_class.sv"
// `include "constraint_outside_class.sv"
// `include "constraint_inheritance.sv"
// `include "constraint_error_scenario.sv"
// `include "constraint_inside_class_02.sv"
// `include "pre_post_randomize.sv"
// `include "inline_constraints.sv"
// `include "inline_with_class_constraints.sv"
// `include "unique_constraint.sv"
// `include "
// `include "
// `include "
// `include "