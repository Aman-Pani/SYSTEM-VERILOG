//`include "array_2d_q3_divisible_by_3or7.sv"
//`include "associative_array_exercise01.sv"
//`include "structure03.sv"
`include "structure04.sv"