// `include "handle_assignment.sv"
// `include "shallow_copy.sv"
// `include "deep_copy.sv"
// `include "class_assignment.sv"
// `include "polymorphism_example.sv"
// `include "inheritance_example01.sv"
`include "encapsulation_example.sv"



