// `include "inheritance01.sv
// `include "q01.sv"
// `include "q02.sv"
// `include "q03.sv"
// `include "parameterized_class.sv"
// `include "scope_resolution.sv"
// `include "typedef_classes.sv"
// `include "casting.sv"
// `include "super.sv"
// `include "overriding.sv"
// `include "polymerphism.sv"
// `include "polymerphism_with_super.sv"
// `include "class_assignment.sv"
// `include "shallow_copy.sv"
`include "deep_copy.sv"
