//write a code to design an array in such a way that the array contains all the numbers those are divisible by 3 or 7 and must bounded in range 50 to 500

module top;
  int d_arr1[int];
  int i,j,count=0;
  
  initial begin
    for(i = 50; i<=500;i++)begin
      if (i % 3 == 0 || i % 7 == 0)begin
        d_arr1[count]=i;
        count++;
      end
    end
    for(j = 0; j<count;j++)begin
      $display(" d_arr1[%0d]=\t %0d",j,d_arr1[j]);
    end
  end
endmodule


// output
//  d_arr1[0]=	 51
//  d_arr1[1]=	 54
//  d_arr1[2]=	 56
//  d_arr1[3]=	 57
//  d_arr1[4]=	 60
//  d_arr1[5]=	 63
//  d_arr1[6]=	 66
//  d_arr1[7]=	 69
//  d_arr1[8]=	 70
//  d_arr1[9]=	 72
//  d_arr1[10]=	 75
//  d_arr1[11]=	 77
//  d_arr1[12]=	 78
//  d_arr1[13]=	 81
//  d_arr1[14]=	 84
//  d_arr1[15]=	 87
//  d_arr1[16]=	 90
//  d_arr1[17]=	 91
//  d_arr1[18]=	 93
//  d_arr1[19]=	 96
//  d_arr1[20]=	 98
//  d_arr1[21]=	 99
//  d_arr1[22]=	 102
//  d_arr1[23]=	 105
//  d_arr1[24]=	 108
//  d_arr1[25]=	 111
//  d_arr1[26]=	 112
//  d_arr1[27]=	 114
//  d_arr1[28]=	 117
//  d_arr1[29]=	 119
//  d_arr1[30]=	 120
//  d_arr1[31]=	 123
//  d_arr1[32]=	 126
//  d_arr1[33]=	 129
//  d_arr1[34]=	 132
//  d_arr1[35]=	 133
//  d_arr1[36]=	 135
//  d_arr1[37]=	 138
//  d_arr1[38]=	 140
//  d_arr1[39]=	 141
//  d_arr1[40]=	 144
//  d_arr1[41]=	 147
//  d_arr1[42]=	 150
//  d_arr1[43]=	 153
//  d_arr1[44]=	 154
//  d_arr1[45]=	 156
//  d_arr1[46]=	 159
//  d_arr1[47]=	 161
//  d_arr1[48]=	 162
//  d_arr1[49]=	 165
//  d_arr1[50]=	 168
//  d_arr1[51]=	 171
//  d_arr1[52]=	 174
//  d_arr1[53]=	 175
//  d_arr1[54]=	 177
//  d_arr1[55]=	 180
//  d_arr1[56]=	 182
//  d_arr1[57]=	 183
//  d_arr1[58]=	 186
//  d_arr1[59]=	 189
//  d_arr1[60]=	 192
//  d_arr1[61]=	 195
//  d_arr1[62]=	 196
//  d_arr1[63]=	 198
//  d_arr1[64]=	 201
//  d_arr1[65]=	 203
//  d_arr1[66]=	 204
//  d_arr1[67]=	 207
//  d_arr1[68]=	 210
//  d_arr1[69]=	 213
//  d_arr1[70]=	 216
//  d_arr1[71]=	 217
//  d_arr1[72]=	 219
//  d_arr1[73]=	 222
//  d_arr1[74]=	 224
//  d_arr1[75]=	 225
//  d_arr1[76]=	 228
//  d_arr1[77]=	 231
//  d_arr1[78]=	 234
//  d_arr1[79]=	 237
//  d_arr1[80]=	 238
//  d_arr1[81]=	 240
//  d_arr1[82]=	 243
//  d_arr1[83]=	 245
//  d_arr1[84]=	 246
//  d_arr1[85]=	 249
//  d_arr1[86]=	 252
//  d_arr1[87]=	 255
//  d_arr1[88]=	 258
//  d_arr1[89]=	 259
//  d_arr1[90]=	 261
//  d_arr1[91]=	 264
//  d_arr1[92]=	 266
//  d_arr1[93]=	 267
//  d_arr1[94]=	 270
//  d_arr1[95]=	 273
//  d_arr1[96]=	 276
//  d_arr1[97]=	 279
//  d_arr1[98]=	 280
//  d_arr1[99]=	 282
//  d_arr1[100]=	 285
//  d_arr1[101]=	 287
//  d_arr1[102]=	 288
//  d_arr1[103]=	 291
//  d_arr1[104]=	 294
//  d_arr1[105]=	 297
//  d_arr1[106]=	 300
//  d_arr1[107]=	 301
//  d_arr1[108]=	 303
//  d_arr1[109]=	 306
//  d_arr1[110]=	 308
//  d_arr1[111]=	 309
//  d_arr1[112]=	 312
//  d_arr1[113]=	 315
//  d_arr1[114]=	 318
//  d_arr1[115]=	 321
//  d_arr1[116]=	 322
//  d_arr1[117]=	 324
//  d_arr1[118]=	 327
//  d_arr1[119]=	 329
//  d_arr1[120]=	 330
//  d_arr1[121]=	 333
//  d_arr1[122]=	 336
//  d_arr1[123]=	 339
//  d_arr1[124]=	 342
//  d_arr1[125]=	 343
//  d_arr1[126]=	 345
//  d_arr1[127]=	 348
//  d_arr1[128]=	 350
//  d_arr1[129]=	 351
//  d_arr1[130]=	 354
//  d_arr1[131]=	 357
//  d_arr1[132]=	 360
//  d_arr1[133]=	 363
//  d_arr1[134]=	 364
//  d_arr1[135]=	 366
//  d_arr1[136]=	 369
//  d_arr1[137]=	 371
//  d_arr1[138]=	 372
//  d_arr1[139]=	 375
//  d_arr1[140]=	 378
//  d_arr1[141]=	 381
//  d_arr1[142]=	 384
//  d_arr1[143]=	 385
//  d_arr1[144]=	 387
//  d_arr1[145]=	 390
//  d_arr1[146]=	 392
//  d_arr1[147]=	 393
//  d_arr1[148]=	 396
//  d_arr1[149]=	 399
//  d_arr1[150]=	 402
//  d_arr1[151]=	 405
//  d_arr1[152]=	 406
//  d_arr1[153]=	 408
//  d_arr1[154]=	 411
//  d_arr1[155]=	 413
//  d_arr1[156]=	 414
//  d_arr1[157]=	 417
//  d_arr1[158]=	 420
//  d_arr1[159]=	 423
//  d_arr1[160]=	 426
//  d_arr1[161]=	 427
//  d_arr1[162]=	 429
//  d_arr1[163]=	 432
//  d_arr1[164]=	 434
//  d_arr1[165]=	 435
//  d_arr1[166]=	 438
//  d_arr1[167]=	 441
//  d_arr1[168]=	 444
//  d_arr1[169]=	 447
//  d_arr1[170]=	 448
//  d_arr1[171]=	 450
//  d_arr1[172]=	 453
//  d_arr1[173]=	 455
//  d_arr1[174]=	 456
//  d_arr1[175]=	 459
//  d_arr1[176]=	 462
//  d_arr1[177]=	 465
//  d_arr1[178]=	 468
//  d_arr1[179]=	 469
//  d_arr1[180]=	 471
//  d_arr1[181]=	 474
//  d_arr1[182]=	 476
//  d_arr1[183]=	 477
//  d_arr1[184]=	 480
//  d_arr1[185]=	 483
//  d_arr1[186]=	 486
//  d_arr1[187]=	 489
//  d_arr1[188]=	 490
//  d_arr1[189]=	 492
//  d_arr1[190]=	 495
//  d_arr1[191]=	 497
//  d_arr1[192]=	 498