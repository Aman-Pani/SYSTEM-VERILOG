class common;
  static mailbox gen2bfm = new();
  static mailbox mon_in2scb = new();
  static mailbox mon_out2scb = new();
  static mailbox mon_in2cov = new();
  static virtual adder_intf vif;
endclass