// https://www.edaplayground.com/x/YG3N

// virtual methods example
// https://www.edaplayground.com/x/4c_p

// pure virtual mehod
// https://www.edaplayground.com/x/62G8

// polymorphism
// https://www.edaplayground.com/x/2Nsi

// abstract class
// https://www.edaplayground.com/x/5K2y
// https://www.edaplayground.com/x/4wqc