// `include "semaphore_01.sv"
// `include "semaphore_02.sv"
`include "semaphore_03_multipleKey.sv"
// `include "
// `include "
// `include "
// `include "
// `include "
// `include "