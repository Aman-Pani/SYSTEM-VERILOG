`include "adder_intf.sv"
`include "common.sv"
`include "adder_tx.sv"
`include "adder_cov.sv"
`include "adder_scb.sv"
`include "adder_mon_out.sv"
`include "adder_mon_in.sv"
`include "adder_gen.sv"
`include "adder_bfm.sv"
`include "adder_agent.sv"
`include "adder_env.sv"
`include "adder_test.sv"
`include "top.sv"