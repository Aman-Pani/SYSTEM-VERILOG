// Code your design here
//module nand_(input a,b,output c);
//  assign c=~(a & b);
//endmodule
module nand_ (
  input a,b
  output c
);
  //assign c=~(a&b);
  assign c=~(a&b);
endmodule