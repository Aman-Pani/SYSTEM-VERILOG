// d12 
// https://www.edaplayground.com/x/LS3R



// virtual_class_basic
// https://www.edaplayground.com/x/5K2y

