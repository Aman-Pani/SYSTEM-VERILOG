// `include "q01_deep_copy_practice.sv"
// `include "q02_method_override.sv"
// `include "q03_method_override_02.sv"
`include "q04.sv"
// `include "virtual_class_basic.sv"
// `include "dynamic_casting.sv"
// `include "extern_method.sv"
// `include "abstract_class.sv"
// `include "mail_box.sv"