// `include "q01.sv"
// `include "q02.sv"
// `include "q03.sv"
// `include "fork_join.sv"
// `include "fork_join_any.sv"
// `include "fork_join_none.sv"
// `include "fork_join_any_waitFork.sv"
// `include "disable_fork.sv"
// `include "disable_fork_example01.sv"
`include "disable_fork_example02.sv"