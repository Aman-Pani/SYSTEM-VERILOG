// `include "practice01_typedef.sv"
// `include "practice02_string.sv"
// `include "practice03_string.sv"
// `include "class01_example.sv"
// `include "class02_example.sv"
// `include "class03_example_thisPointer_wo.sv"
// `include "class04_example_thisPointer_w.sv"
// `include "class05_example_constructor.sv"
// `include "class06_example_thisPointer_w_02.sv"
// `include "class07_example_staticVariable.sv"
// `include "class08_example_staticVariable.sv"
// `include "class09_example_staticVariable.sv"
`include "class10_example_staticVariable.sv"