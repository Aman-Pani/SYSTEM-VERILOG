class common;
  static mailbox gen2bfm = new();
  static virtual adder_intf vif;
endclass