// d14 :	https://www.edaplayground.com/x/kzFP